// For loop - For loop is use to execute the statements again and agains .When the condition ofr for loop 
//          will not true , it will get terminate and the user will come out from the loop .
//  Syntax - // declaring the data type to the variable 
//              assign the value to the variable 
//              initial begin 
//              for ([initialization]; [condition]; [modifier])
//               begin 
//               Statements;
//               end
//               end// 
//               
// Example - 
//
module for_code;

        



